---------------------------------------------------------------------------------------------------------------------
	-- COMPANY: TECHNICAL UNIVERSITY OF CRETE
	-- ENGINEER: NICK KYPARISSAS
	-- 
	-- CREATE DATE: 14 JUNE 2015 
	-- DESIGN NAME: 
	-- MODULE NAME: CELLULAR_AUTOMATON_MODULE - BEHAVIORAL
	-- TARGET DEVISES: SYNTHESIZABLE, A VARIATION HAS BEEN TESTED ON NEXYS 4.
	--
	-- DESCRIPTION: THIS MODULE LOADS AN EXANDING CELLULAR AUTOMATON (CA) FROM MEMORY MODULE NO. 1, 
	-- ACTS ON IT ACCORDING TO THE CA'S RULES AND STORES THE RESULT IN MEMORY MODULE NO. 2. 
	-- THEN IT EXCHANGES THE MEMORY MODULES, READS FROM MEMORY MODULE NO. 2 AND WRITES IN MEMORY MODULE NO. 1.
	-- DUE TO LIMITED MEMORY SIZE, I HAD TO AVOID HAVING DYING CELLS (BECAUSE THEN YOU NEED MORE MEMORY TO 
	-- STORE A 3RD FRAME WITHOUT ANY CELLS ON IT), SO THIS MODULE IMPLEMENTS A FOREVER EXPANDING CA.
	--
	-- IMPLEMENTED FOR XILINX UNIVERSITY PROGRAM'S "OPEN HARDWARE 2015" COMPETITION.
---------------------------------------------------------------------------------------------------------------------


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CELLULAR_AUTOMATON_MODULE IS
	GENERIC(
		GRID_SIZE_X  		:  INTEGER := 100; -- USUALLY FITS INTO A SCREEN RESOLUTION, A MEMORY OR A SUBDIVISION OF THOSE.
		GRID_SIZE_Y  		:  INTEGER := 100;
		NEIGHBORHOOD_SIZE 	: INTEGER := 3 -- MOORE NEIGHBORHOOD SIZE: USE "3" FOR THE CLASSIC 3X3 MOORE NEIGHBORHOOD.
	);
	PORT ( DATA_IN          : IN STD_LOGIC_VECTOR (7 DOWNTO 0); -- DATA SIZE, HERE: A BYTE.
		EN               	: IN STD_LOGIC; -- WHEN EN COMES, IT EXCHANGES BETWEEN THE TWO MEMORY MODULES.
		RST              	: IN STD_LOGIC;
		CLOCK            	: IN STD_LOGIC;
		WEN              	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		SEL              	: OUT STD_LOGIC;
		ADDRESS          	: OUT STD_LOGIC_VECTOR (13 DOWNTO 0); -- IT NEEDS TO FIT THE GRID AND THE MEMORY. 
	DATA_OUT         : OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
END CELLULAR_AUTOMATON_MODULE;

ARCHITECTURE BEHAVIORAL OF CELLULAR_AUTOMATON_MODULE IS
	
	TYPE STATE IS (RESET, READ, STORE, CALCULATE_CA_INITIALIZATION, CALCULATE_CA, WRITE, CALCULATE_NEXT_CELL, WAIT_EN, EX_MEM);
	SIGNAL Y 				: STATE;
	SIGNAL CURRENT_CELL_X 	: STD_LOGIC_VECTOR(6 DOWNTO 0); -- IT NEEDS TO FIT THE GRID_SIZE_X'S MAXIMUM VALUE. SET IT AS THE CENTRAL CELL'S X DIMENSION OF THE FIRST FULL NEIGHBORHOOD OF YOUR GRID. FOR EXAMPLE, FOR A 7X7 GRID, IT'S VALUE WOULD BE 3.
	SIGNAL CURRENT_CELL_Y 	: STD_LOGIC_VECTOR(13 DOWNTO 0); -- IT NEEDS TO FIT THE (GRID_SIZE_X * GRID_SIZE_Y)'S MAXIMUM VALUE.
	SIGNAL GRID_X 			: STD_LOGIC_VECTOR(6 DOWNTO 0); -- DIMENSIONS OF THE CELL TO BE READ OR WRITTEN. AT FIRST, IT HAS TO BE THE FIRST CELL OF THE NEIGHBORHOOD. 
	SIGNAL GRID_Y 			: STD_LOGIC_VECTOR(13 DOWNTO 0); 
	SIGNAL COUNTER 			: STD_LOGIC_VECTOR(3 DOWNTO 0); -- IT NEEDS TO FIT NEIGHBORHOOD_SIZE^2.
	SIGNAL SEL_SIG 			: STD_LOGIC;

BEGIN 
	
	CA_RULES: PROCESS 
		BEGIN
		
		WAIT UNTIL CLOCK'EVENT AND CLOCK = '1';
		
		IF ( RST = '1' ) THEN  
		Y <= RESET;    
		ELSE
			CASE Y IS 
				WHEN RESET =>
					-- OUTPUTS:
					SEL_SIG <= '0'; -- SELECT THE FIRST RAM MODULE.
					WEN <= "0"; -- DO NOT WRITE ANYTHING.
					-- THE OTHER OUTPUTS' VALUES ARE IRRELEVANT HERE.
					-- SIGNALS:
					CURRENT_CELL_X <= "0000001"; -- THE CENTRAL CELL'S X DIMENSION OF THE FIRST FULL NEIGHBORHOOD, HERE: 1X1.
					CURRENT_CELL_Y <= "00000001100100"; -- CURRENT_CELL_Y IS COMPUTED AS: CURRENT ROW'S NUMBER * GRID_SIZE_X.  
					GRID_X <= (OTHERS => '0'); -- INITIATE ADDRESS 0, FIRST CELL OF THE GRID - FIRST CELL OF THE FIRST NEIGHBORHOOD.
					GRID_Y <= (OTHERS => '0');
					COUNTER <= (OTHERS => '0');
					-- NEXT STATE:
					Y <= READ;
				WHEN STORE =>
					IF (GRID_X = CURRENT_CELL_X + NEIGHBORHOOD_SIZE/2) AND (GRID_Y = CURRENT_CELL_Y + GRID_SIZE_X*NEIGHBORHOOD_SIZE/2) THEN --IF THE FINAL CELL OF THE NEIGHBORHOOD.
						GRID_X <= CURRENT_CELL_X;
						GRID_Y <= CURRENT_CELL_Y;
						Y <= CALCULATE_CA_INITIALIZATION;
					ELSE -- CALCULATE NEXT ADDRESS.
						IF (GRID_X = CURRENT_CELL_X + NEIGHBORHOOD_SIZE/2) THEN 
							GRID_X <= CURRENT_CELL_X - NEIGHBORHOOD_SIZE/2; -- THE FIRST CELL OF THE NEXT ROW OF THE NEIGHBORHOOD.
							GRID_Y <= GRID_Y + GRID_SIZE_X;
						ELSE
							GRID_X <= GRID_X + 1;
						END IF;
						Y <= READ;
					END IF;
					-- CHECK THE MOORE NEIGHBORHOOD (NOT THE EXTENDED ONE, BUT THE NORMAL 3X3 NEIGHBORHOOD).
					IF (GRID_Y > CURRENT_CELL_Y - 2*GRID_SIZE_X) AND (GRID_Y < CURRENT_CELL_Y + 2*GRID_SIZE_X) AND (GRID_X > CURRENT_CELL_X - 2) AND (GRID_X < CURRENT_CELL_X + 2) THEN
						IF (DATA_IN /= "00000000") THEN --IF WE HAVE DATA IN THE NEIGHBORHOOD.
							COUNTER <= COUNTER + 1;
						END IF;
					END IF;
					-- STORE THE APPROPRIATE COUNTER VALUES.
					IF (GRID_X /= CURRENT_CELL_X) AND (GRID_Y /= CURRENT_CELL_Y) THEN -- IF WE ARE NOT READING THE CURRENT CELL.
						IF (DATA_IN /= "00000000") THEN -- IF WE HAVE DATA IN THE EXTENDED NEIGHBORHOOD. YOU CAN INCREASE DIFFERENT COUNTERS FOR DIFFERENT TYPES OF DATA! 
							COUNTER <= COUNTER + 1;
						END IF; 
					END IF; 
				WHEN READ =>   -- THE ADDRESSES HERE HAVE BEEN SET. IN THE NEXT CYCLE, THE DATA WILL HAVE BEEN SET ON THE DATA BUS.
					Y <= STORE;                     
				WHEN CALCULATE_CA_INITIALIZATION => --THE ADDRESSES HERE HAVE BEEN SET. IN THE NEXT CYCLE, THE DATA WILL HAVE BEEN SET ON THE DATA BUS.
					Y <= CALCULATE_CA;    
				WHEN CALCULATE_CA =>
					IF (COUNTER > 3) THEN -- IF THE RULES APPLY, FOR EXAMPLE HERE: COUNTER > 3
						DATA_OUT <= "10101010"; -- WRITE WHAT THE RULES SAY.
					ELSE 
						DATA_OUT <= DATA_IN;      
					END IF;
					WEN <= "1";
					Y <= WRITE;
				WHEN WRITE => -- IF WE ARE IN THE END OF THE FRAME.
					IF ((CURRENT_CELL_X = GRID_SIZE_X - NEIGHBORHOOD_SIZE/2) AND (CURRENT_CELL_Y = GRID_SIZE_X*(GRID_SIZE_Y-1))) THEN -- FINAL CELL
						Y <= WAIT_EN; -- THIS "WAIT" STATE HAS BEEN SET IN CASE YOU WANT TO CONTROL THE CA'S SPEED. IF YOU DON'T WANT THAT, JUMP TO "EX_MEM".  
					ELSE
						Y <= CALCULATE_NEXT_CELL;
					END IF; 
					WEN <= "0";
				WHEN CALCULATE_NEXT_CELL =>
					IF (CURRENT_CELL_X = GRID_SIZE_X - NEIGHBORHOOD_SIZE/2) THEN
						CURRENT_CELL_X <= "0000001"; -- THE CENTRAL CELL'S X DIMENSION OF THE FIRST FULL NEIGHBORHOOD, HERE: 1X1.
						CURRENT_CELL_Y <= CURRENT_CELL_Y + GRID_SIZE_X; --CHANGE LINE
						GRID_X <= (OTHERS => '0'); -- INITIATE ADDRESS POINTING AT THE FIRST CELL OF THE NEXT NEIGHBORHOOD.
						GRID_Y <= STD_LOGIC_VECTOR(TO_UNSIGNED(NEIGHBORHOOD_SIZE/2, GRID_Y'LENGTH));
					ELSE
						CURRENT_CELL_X <= CURRENT_CELL_X + 1;
						GRID_X <= CURRENT_CELL_X - NEIGHBORHOOD_SIZE/2 -1; -- INITIATE ADDRESS POINTING AT THE FIRST CELL OF THE NEXT NEIGHBORHOOD.
						GRID_Y <= CURRENT_CELL_Y - GRID_SIZE_X*NEIGHBORHOOD_SIZE/2;
					END IF;
					COUNTER <= (OTHERS => '0');
					Y <= READ;
				WHEN WAIT_EN => -- THIS "WAIT" STATE HAS BEEN SET IN CASE YOU WANT TO CONTROL THE CA'S SPEED.
					IF (EN = '1') THEN
						Y <= EX_MEM;
					ELSE
						Y <= Y;
					END IF;
				WHEN EX_MEM =>
					SEL_SIG <= NOT SEL_SIG; -- NEXT FRAME, EXCHANGE MEMORIES. 
					-- SIGNALS:
					CURRENT_CELL_X <= "0000001"; -- THE CENTRAL CELL'S X DIMENSION OF THE FIRST FULL NEIGHBORHOOD, HERE: 1X1.
					CURRENT_CELL_Y <= "00000001100100"; -- CURRENT_CELL_Y IS COMPUTED AS: CURRENT ROW'S NUMBER * GRID_SIZE_X.  
					GRID_X <= (OTHERS => '0'); -- INITIATE ADDRESS 0, FIRST CELL OF THE GRID - FIRST CELL OF THE FIRST NEIGHBORHOOD
					GRID_Y <= (OTHERS => '0');
					COUNTER <= (OTHERS => '0');
					Y <= READ;
			END CASE;  
		END IF;                    
	END PROCESS CA_RULES;
	
	ADDRESS <= GRID_X + GRID_Y;
	SEL <= SEL_SIG;

END BEHAVIORAL;